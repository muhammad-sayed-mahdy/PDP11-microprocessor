LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

--Control Store
ENTITY rom IS
	GENERIC ( n : integer := 21);
	PORT(
		address : IN  std_logic_vector(5 DOWNTO 0);
		dataout : OUT std_logic_vector(n-1 DOWNTO 0));
END ENTITY rom;

ARCHITECTURE rom_arch OF rom IS

	TYPE rom_type IS ARRAY(0 TO 63) OF std_logic_vector(n-1 DOWNTO 0);
	SIGNAL rom : rom_type := (
		"110101000101101010101",
		"000100010000000100000",
		"000100001000000100000",
		"000010010000001000001",
		"001000010100000010000",
		"000111010001101010101",
		"000010001000001000001",
		"000010001110000000000",
		"001010011001100001100",
		"110111010001100011000",
		"000000001110100000000",
		"000000001100010000010",
		"010000010100001000001",
		"001111000101101010101",
		"001000010100001000000",
		"010001001100100000000",
		"001000001000000010000",
		"010010001000000010000",
		"010011010001100000000",
		"000010001100001000001",
		"010101010101101010101",
		"000000001110100000000",
		"000000001110101000001",
		"011001001100100000000",
		"010000001000001000001",
		"011011001000000010000",
		"001000001000001000000",
		"011100010101100000000",
		"000000001100001000001",
		"011110001100100000000",
		"011111001000000100000",
		"100000100001100011000",
		"100001001111001000000",
		"100010000100010000010",
		"000000011000100000000",
		"100101001111000000000",
		"010110010101100011000",
		"000000001000100000000",
		"100111100001100011000",
		"101001001111001000010",
		"110001100101100011100",
		"101010000100010000000",
		"101011100001100011000",
		"111111001111001000010",
		"101101001111000000000",
		"101110001000100000000",
		"101111100001101010101",
		"110000001111000000000",
		"000000001011100000000",
		"110010001100000010000",
		"110011000101100000000",
		"000000001100100000000",
		"010111000101101010101",
		"110110001100100000000",
		"000000001001000000000",
		"000010001110001000001",
		"011101000101101010101",
		"100011100001101010101",
		"101100100001101010101",
		"100110011100010000000",
		"000000011010100000000",
		"000000000000000000000",
		"000000011000010000010",
		"111111000000000000000"
	);
	BEGIN
		dataout <= rom(to_integer(unsigned(address)));
END rom_arch;
